package soc_pkg ; 



  import uvm_pkg::*;
`include "uvm_macros.svh"


// import uart_pkg::*;
// import wb_pkg::*;

`include "soc_ref_env.sv.sv"
`include "soc_scb.sv"
`include "soc_ref_model.sv.sv"



endpackage